`timescale 1ns / 1ps

module fa_fs_tb;
reg a,b,cin;
wire s,ca,di,bo;

fa_fs_mux dut(a,b,cin,s,ca,di,bo);
initial
    begin
    a=0;b=0;cin=0;
    #10 a=0;b=0;cin=1;
    #10 a=0;b=1;cin=0;
    #10 a=0;b=1;cin=1;
    #10 a=1;b=0;cin=0;
    #10 a=1;b=0;cin=1;
    #10 a=1;b=1;cin=0;
    #10 a=1;b=1;cin=1;
    #10 $finish;
    
    
    end
endmodule